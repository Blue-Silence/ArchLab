`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Create Date: 2023/02/07 15:21:49
//////////////////////////////////////////////////////////////////////////////////


module Decoder(input [3:0] i , output [6:0] o);

    assign o = (i==0) ? 7'b1000000 :
               (i==1) ? 7'b1111001 : 
               (i==2) ? 7'b0100100 :
               (i==3) ? 7'b0110000 :
               (i==4) ? 7'b0011001 :
               (i==5) ? 7'b0010010 :
               (i==6) ? 7'b0000010 :
               (i==7) ? 7'b1111000 :
               (i==8) ? 7'b0000000 :
               (i==9) ? 7'b0010000 :
               (i==10) ? 7'b0001000 :
               (i==11) ? 7'b0000011 :
               (i==12) ? 7'b1000110 :
               (i==13) ? 7'b0100001 :
               (i==14) ? 7'b0000110 :
               (i==15) ? 7'b0001110 :
               7'bx ;
               
endmodule
